

`define m_bits       4   
`define id_bits      6
`define slave_id_bits 7
`define addr_bits   44
`define len_bits     8
`define data_bits  128
`define strb_bits    (`data_bits/8)
`define size_bits    3
`define burst_bits   2
`define lock_bits    1
`define cache_bits   4
`define prot_bits    3
`define resp_bits    4
`define ruser_bits   7
`define wuser_bits   9
`define snoop_bits   3
